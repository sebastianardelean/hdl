//----------------------------------------------
// Design Name:  
// File Name: 
// Function: 
// Version | Changes | Author
//----------------------------------------------
