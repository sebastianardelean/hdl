`ifndef __DEFS_SVH__
 `define __DEFS_SVH__

`timescale 1ns/1ps


`endif // __DEFS_SVH__
