`ifndef __DEFS_SVH__
 `define __DEFS_SVH__




`endif // __DEFS_SVH__
